library verilog;
use verilog.vl_types.all;
entity ID_EX_Reg is
    port(
        RegWriteD       : in     vl_logic;
        ResultSrcD      : in     vl_logic_vector(2 downto 0);
        MemWriteD       : in     vl_logic;
        MemReadD        : in     vl_logic;
        JumpD           : in     vl_logic;
        JumpTypeD       : in     vl_logic;
        BranchD         : in     vl_logic;
        BranchTypeD     : in     vl_logic_vector(2 downto 0);
        ALUControlD     : in     vl_logic_vector(2 downto 0);
        ALUSrcD         : in     vl_logic;
        SLTControlD     : in     vl_logic_vector(1 downto 0);
        StrobeD         : in     vl_logic_vector(2 downto 0);
        mretD           : in     vl_logic;
        csrOpD          : in     vl_logic_vector(1 downto 0);
        CUexceptionD    : in     vl_logic;
        CUexceptionTypeD: in     vl_logic_vector(3 downto 0);
        RD1D            : in     vl_logic_vector(31 downto 0);
        RD2D            : in     vl_logic_vector(31 downto 0);
        InstrD          : in     vl_logic_vector(31 downto 0);
        PCD             : in     vl_logic_vector(31 downto 0);
        Rs1D            : in     vl_logic_vector(4 downto 0);
        Rs2D            : in     vl_logic_vector(4 downto 0);
        RdD             : in     vl_logic_vector(4 downto 0);
        ExtImmD         : in     vl_logic_vector(31 downto 0);
        PCPlus4D        : in     vl_logic_vector(31 downto 0);
        rst             : in     vl_logic;
        clk             : in     vl_logic;
        EN              : in     vl_logic;
        FLUSH           : in     vl_logic;
        RegWriteE       : out    vl_logic;
        ResultSrcE      : out    vl_logic_vector(2 downto 0);
        MemWriteE       : out    vl_logic;
        MemReadE        : out    vl_logic;
        JumpE           : out    vl_logic;
        JumpTypeE       : out    vl_logic;
        BranchE         : out    vl_logic;
        BranchTypeE     : out    vl_logic_vector(2 downto 0);
        ALUControlE     : out    vl_logic_vector(2 downto 0);
        ALUSrcE         : out    vl_logic;
        SLTControlE     : out    vl_logic_vector(1 downto 0);
        StrobeE         : out    vl_logic_vector(2 downto 0);
        mretE           : out    vl_logic;
        csrOpE          : out    vl_logic_vector(1 downto 0);
        CUexceptionE    : out    vl_logic;
        CUexceptionTypeE: out    vl_logic_vector(3 downto 0);
        RD1E            : out    vl_logic_vector(31 downto 0);
        RD2E            : out    vl_logic_vector(31 downto 0);
        Rs1E            : out    vl_logic_vector(4 downto 0);
        Rs2E            : out    vl_logic_vector(4 downto 0);
        RdE             : out    vl_logic_vector(4 downto 0);
        ExtImmE         : out    vl_logic_vector(31 downto 0);
        InstrE          : out    vl_logic_vector(31 downto 0);
        PCE             : out    vl_logic_vector(31 downto 0);
        PCPlus4E        : out    vl_logic_vector(31 downto 0)
    );
end ID_EX_Reg;
