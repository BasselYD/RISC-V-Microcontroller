library verilog;
use verilog.vl_types.all;
entity Test_tb is
end Test_tb;
